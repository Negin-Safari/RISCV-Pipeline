module inst_mem (adr, d_out);
  input [64:0] adr;
  output [31:0] d_out;
  
  reg [7:0] mem[0:65535];
  
  initial
  begin
    //         add    R8, R0, R0 0
    //         addi   R10,  R0, 20 4
    //         ld     R2, 1000(R8) 8
    //         add    R3, R0, R8    12
    // Loop:   beq    R8,  R10, END_LOOP 16   
    //         add    R13, R8, R8      20     /////
    //         add    R13, R13, R13     24    ////
    //         add    R13, R13, R13     28
    //         ld     R7, 1000(R13)     32      ///
    //         slt    R11, R7, R2       36 
    //         beq    R0, R11, END_IF   40    ////////////////
    //    	    add    R2, R0, R7        44  //////
    //         add    R3, R0, R8        48
    // END_IF: addi   R8, R8, 1         52
    //         J      LOOP              56   ////(beq)
    // END_LOOP: sd, R2, 2000(R0)       60
    //           sd, R3, 2004(R0)       64
    ///////////////// // 
    //            jal  X1, TEST         68
    //  RETURTN:  sll R17,R3,R2         72
    //            srl R18,R3,R2         76
    
    //  TEST:     sub R9,R3,R2          120
    //            or R12,R3,R2          124
    //            and R14,R3,R2         128
    //            slti R15,R2,20        132
    //            jalr R16 RETURN(R2)   136

    
//   {mem[3], mem[2], mem[1], mem[0]}     = {7'd0, 5'd0, 5'd0,3'd0, 5'd8,7'b0110011};   
//   {mem[7], mem[6], mem[5], mem[4]}     = {12'd20, 5'd0,3'd0, 5'd10, 7'b0010011};               
//   {mem[11], mem[10], mem[9], mem[8]}   = {12'd1000, 5'd8, 3'd3,5'd2,7'b0000011};                
//   {mem[15], mem[14], mem[13], mem[12]} = {7'd0, 5'd8, 5'd0, 3'd0, 5'd3,7'b0110011};           
//   {mem[19], mem[18], mem[17], mem[16]} = {1'd0,6'd1,5'd10,5'd8,3'd0,4'd6,1'd0,7'b1100011};  ////
//   {mem[23], mem[22], mem[21], mem[20]} = {7'd0, 5'd8, 5'd8,3'd0,5'd13,7'b0110011};              
//   {mem[27], mem[26], mem[25], mem[24]} = {7'd0, 5'd13, 5'd13,3'd0,5'd13,7'b0110011}; 
//   {mem[31], mem[30], mem[29], mem[28]} = {7'd0, 5'd13, 5'd13,3'd0,5'd13,7'b0110011};           
//   {mem[35], mem[34], mem[33], mem[32]} = {12'd1000, 5'd13, 3'd3,5'd7,7'b0000011};
//   {mem[39], mem[38], mem[37], mem[36]} = {7'd0, 5'd2, 5'd7, 3'd2, 5'd11, 7'b0110011}; 
//   {mem[43], mem[42], mem[41], mem[40]} = {1'd0, 6'd0, 5'd11, 5'd0, 3'd0, 4'd6, 1'd0,7'b1100011}; 
//   {mem[47], mem[46], mem[45], mem[44]} = {7'd0, 5'd7, 5'd0,3'd0, 5'd2,7'b0110011};
//   {mem[51], mem[50], mem[49], mem[48]} = {7'd0, 5'd8, 5'd0,3'd0, 5'd3,7'b0110011};
//   {mem[55], mem[54], mem[53], mem[52]} = {12'd1, 5'd8,3'd0, 5'd8, 7'b0010011}; 
//   {mem[59], mem[58], mem[57], mem[56]} = {1'd1, 6'd62,5'd0,5'd0,3'd0,4'd12,1'd1,7'b1100011}; ////
//   {mem[63], mem[62], mem[61], mem[60]} = {7'd62, 5'd2, 5'd0, 3'd7, 5'd16, 7'b0100011};
//   {mem[67], mem[66], mem[65], mem[64]} = {7'd62, 5'd3, 5'd0, 3'd7, 5'd24, 7'b0100011}; 
     $readmemb( "INST.mem", mem ); 
//// srl,sll,jal,jalr,slti,lw,sw
//   {mem[71], mem[70], mem[69], mem[68]} = {1'd0,10'd26,1'd0,8'd0,5'd1,7'b1101111};	 //dorost shoo
//   {mem[75], mem[74], mem[73], mem[72]} = {7'd0,5'd2,5'd3,3'd1,5'd17,7'b0110011};
//   {mem[79], mem[78], mem[77], mem[76]} = {7'd0,5'd2,5'd3,3'd5,5'd18,7'b0110011};

//   {mem[123], mem[122], mem[121], mem[120]} = {7'd32,5'd2,5'd3,3'd0,5'd9,7'b0110011};
//   {mem[127], mem[126], mem[125], mem[124]} = {7'd0,5'd2,5'd3,3'd6,5'd12,7'b0110011};
//   {mem[131], mem[130], mem[129], mem[128]} = {7'd0,5'd2,5'd3,3'd7,5'd14,7'b0110011};
//   {mem[135], mem[134], mem[133], mem[132]} = {12'd20,5'd2,3'd2,5'd15,7'b0010011};
//   {mem[139], mem[138], mem[137], mem[136]} = {-12'd35,5'd2,3'd0,5'd16,7'b1100111};
    
  end
  
  assign d_out = {mem[adr[15:0]+3], mem[adr[15:0]+2], mem[adr[15:0]+1], mem[adr[15:0]]};
  
endmodule
